SQRT_inst : SQRT PORT MAP (
		clk	 => clk_sig,
		radical	 => radical_sig,
		q	 => q_sig,
		remainder	 => remainder_sig
	);
